class seqr extends uvm_sequencer#(seqt);
`uvm_component_utils(seqr)

`compnew

endclass
