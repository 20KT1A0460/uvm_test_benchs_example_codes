     interface interf1();  //single interface to both mux and decoder
     logic [3:0] a,b,c,d,y; //mux ports
     logic s1,s2;  
     logic f,g,y1,y2,y3,y4; //decoder ports
     endinterface




