interface interf();
logic [3:0]a,b,sum;
logic cin,carry;
endinterface

interface interf2();
logic [3:0]a,b,sum;
logic cin,carry;
endinterface
